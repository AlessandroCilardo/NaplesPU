//        Copyright 2019 NaplesPU
//   
//   	 
//   Redistribution and use in source and binary forms, with or without modification,
//   are permitted provided that the following conditions are met:
//   
//   1. Redistributions of source code must retain the above copyright notice,
//      this list of conditions and the following disclaimer.
//   
//   2. Redistributions in binary form must reproduce the above copyright notice,
//      this list of conditions and the following disclaimer in the documentation
//      and/or other materials provided with the distribution.
//   
//   3. Neither the name of the copyright holder nor the names of its contributors
//      may be used to endorse or promote products derived from this software
//      without specific prior written permission.
//   
//      
//   THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//   ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//   WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
//   IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
//   INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
//   BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
//   DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
//   LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE
//   OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED
//   OF THE POSSIBILITY OF SUCH DAMAGE.

`timescale 1ns / 1ps
module priority_encoder_npu #(
        parameter INPUT_WIDTH   = 4,
        parameter MAX_PRIORITY  = "LSB"
    )(
        input   logic   [INPUT_WIDTH            - 1 : 0]    decode,
        output  logic   [$clog2(INPUT_WIDTH)    - 1 : 0]    encode,
        output  logic                                       valid
    );

    generate
        always_comb begin
            encode = 0;
            if (MAX_PRIORITY == "LSB") begin
                for (int i = INPUT_WIDTH - 1; i >= 0; i--)
                    if (decode[i] == 1)
                        encode = i[$clog2(INPUT_WIDTH)  - 1 : 0];
            end else begin
                for (int i = 0; i < INPUT_WIDTH; i++)
                    if (decode[i] == 1)
                        encode = i[$clog2(INPUT_WIDTH)  - 1 : 0];
            end
        end
    endgenerate

    assign valid = |decode;

endmodule
