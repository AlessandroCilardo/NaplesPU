//        Copyright 2019 NaplesPU
//   
//   	 
//   Redistribution and use in source and binary forms, with or without modification,
//   are permitted provided that the following conditions are met:
//   
//   1. Redistributions of source code must retain the above copyright notice,
//      this list of conditions and the following disclaimer.
//   
//   2. Redistributions in binary form must reproduce the above copyright notice,
//      this list of conditions and the following disclaimer in the documentation
//      and/or other materials provided with the distribution.
//   
//   3. Neither the name of the copyright holder nor the names of its contributors
//      may be used to endorse or promote products derived from this software
//      without specific prior written permission.
//   
//      
//   THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
//   ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
//   WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
//   IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
//   INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
//   BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
//   DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF
//   LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE
//   OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED
//   OF THE POSSIBILITY OF SUCH DAMAGE.

`timescale 1ns / 1ps

module grant_hold_round_robin_arbiter
    #(parameter SIZE = 4)

    (input                    clk,
    input                     reset,
    input[SIZE - 1:0]         requests,
    input[SIZE - 1:0]         hold_in,
    output logic[SIZE - 1:0]  decision_oh);

	logic anyhold;
	logic [SIZE - 1:0] grant_arb,last,hold;

	round_robin_arbiter #(
		.SIZE(SIZE)
	)
	u_round_robin_arbiter (
		.clk         ( clk       ),
		.reset       ( reset     ),
		.en          ( 1'b0      ), 
		//.en          ('{default:'0}),
		.requests    ( requests   ),
		.decision_oh ( grant_arb )
	);
	
	assign decision_oh = anyhold ? hold : grant_arb ;
	assign hold = last & hold_in;
	assign anyhold = | hold;
	
	always_ff @(posedge clk, posedge reset) begin
	    if (reset) 
	    	last <= 0;
	    else
	    	last <= decision_oh;   
	end

endmodule

